module _32_bit_and(out,a,b);

input [31:0]a;
input [31:0]b;
output [31:0]out;

and a1(out[0],a[0],b[0]);
and a2(out[1],a[1],b[1]);
and a3(out[2],a[2],b[2]);
and a4(out[3],a[3],b[3]);
and a5(out[4],a[4],b[4]);
and a6(out[5],a[5],b[5]);
and a7(out[6],a[6],b[6]);
and a8(out[7],a[7],b[7]);
and a9(out[8],a[8],b[8]);
and a10(out[9],a[9],b[9]);
and a11(out[10],a[10],b[10]);
and a12(out[11],a[11],b[11]);
and a13(out[12],a[12],b[12]);
and a14(out[13],a[13],b[13]);
and a15(out[14],a[14],b[14]);
and a16(out[15],a[15],b[15]);
and a17(out[16],a[16],b[16]);
and a18(out[17],a[17],b[17]);
and a19(out[18],a[18],b[18]);
and a20(out[19],a[19],b[19]);
and a21(out[20],a[20],b[20]);
and a22(out[21],a[21],b[21]);
and a23(out[22],a[22],b[22]);
and a24(out[23],a[23],b[23]);
and a25(out[24],a[24],b[24]);
and a26(out[25],a[25],b[25]);
and a27(out[26],a[26],b[26]);
and a28(out[27],a[27],b[27]);
and a29(out[28],a[28],b[28]);
and a30(out[29],a[29],b[29]);
and a31(out[30],a[30],b[30]);
and a32(out[31],a[31],b[31]);

endmodule