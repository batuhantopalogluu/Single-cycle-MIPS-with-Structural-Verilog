module shift_right_logic(a,b,out);
	
input[31:0] a;
input[31:0] b;
output[31:0] out;

wire[31:0] tempResult0,tempResult1,tempResult2,tempResult3,temp_out;
wire overflow;
wire not_overflow;


_2_1_mux_v2 mux_layer0_1(a[0],a[1],b[0],tempResult0[0]);
_2_1_mux_v2 mux_layer0_2(a[1],a[2],b[0],tempResult0[1]);
_2_1_mux_v2 mux_layer0_3(a[2],a[3],b[0],tempResult0[2]);
_2_1_mux_v2 mux_layer0_4(a[3],a[4],b[0],tempResult0[3]);
_2_1_mux_v2 mux_layer0_5(a[4],a[5],b[0],tempResult0[4]);
_2_1_mux_v2 mux_layer0_6(a[5],a[6],b[0],tempResult0[5]);
_2_1_mux_v2 mux_layer0_7(a[6],a[7],b[0],tempResult0[6]);
_2_1_mux_v2 mux_layer0_8(a[7],a[8],b[0],tempResult0[7]);
_2_1_mux_v2 mux_layer0_9(a[8],a[9],b[0],tempResult0[8]);
_2_1_mux_v2 mux_layer0_10(a[9],a[10],b[0],tempResult0[9]);
_2_1_mux_v2 mux_layer0_11(a[10],a[11],b[0],tempResult0[10]);
_2_1_mux_v2 mux_layer0_12(a[11],a[12],b[0],tempResult0[11]);
_2_1_mux_v2 mux_layer0_13(a[12],a[13],b[0],tempResult0[12]);
_2_1_mux_v2 mux_layer0_14(a[13],a[14],b[0],tempResult0[13]);
_2_1_mux_v2 mux_layer0_15(a[14],a[15],b[0],tempResult0[14]);
_2_1_mux_v2 mux_layer0_16(a[15],a[16],b[0],tempResult0[15]);
_2_1_mux_v2 mux_layer0_17(a[16],a[17],b[0],tempResult0[16]);
_2_1_mux_v2 mux_layer0_18(a[17],a[18],b[0],tempResult0[17]);
_2_1_mux_v2 mux_layer0_19(a[18],a[19],b[0],tempResult0[18]);
_2_1_mux_v2 mux_layer0_20(a[19],a[20],b[0],tempResult0[19]);
_2_1_mux_v2 mux_layer0_21(a[20],a[21],b[0],tempResult0[20]);
_2_1_mux_v2 mux_layer0_22(a[21],a[22],b[0],tempResult0[21]);
_2_1_mux_v2 mux_layer0_23(a[22],a[23],b[0],tempResult0[22]);
_2_1_mux_v2 mux_layer0_24(a[23],a[24],b[0],tempResult0[23]);
_2_1_mux_v2 mux_layer0_25(a[24],a[25],b[0],tempResult0[24]);
_2_1_mux_v2 mux_layer0_26(a[25],a[26],b[0],tempResult0[25]);
_2_1_mux_v2 mux_layer0_27(a[26],a[27],b[0],tempResult0[26]);
_2_1_mux_v2 mux_layer0_28(a[27],a[28],b[0],tempResult0[27]);
_2_1_mux_v2 mux_layer0_29(a[28],a[29],b[0],tempResult0[28]);
_2_1_mux_v2 mux_layer0_30(a[29],a[30],b[0],tempResult0[29]);
_2_1_mux_v2 mux_layer0_31(a[30],a[31],b[0],tempResult0[30]);
_2_1_mux_v2 mux_layer0_32(a[31],1'b0,b[0],tempResult0[31]);

_2_1_mux_v2 mux_layer1_1(tempResult0[0],tempResult0[2],b[1],tempResult1[0]);
_2_1_mux_v2 mux_layer1_2(tempResult0[1],tempResult0[3],b[1],tempResult1[1]);
_2_1_mux_v2 mux_layer1_3(tempResult0[2],tempResult0[4],b[1],tempResult1[2]);
_2_1_mux_v2 mux_layer1_4(tempResult0[3],tempResult0[5],b[1],tempResult1[3]);
_2_1_mux_v2 mux_layer1_5(tempResult0[4],tempResult0[6],b[1],tempResult1[4]);
_2_1_mux_v2 mux_layer1_6(tempResult0[5],tempResult0[7],b[1],tempResult1[5]);
_2_1_mux_v2 mux_layer1_7(tempResult0[6],tempResult0[8],b[1],tempResult1[6]);
_2_1_mux_v2 mux_layer1_8(tempResult0[7],tempResult0[9],b[1],tempResult1[7]);
_2_1_mux_v2 mux_layer1_9(tempResult0[8],tempResult0[10],b[1],tempResult1[8]);
_2_1_mux_v2 mux_layer1_10(tempResult0[9],tempResult0[11],b[1],tempResult1[9]);
_2_1_mux_v2 mux_layer1_11(tempResult0[10],tempResult0[12],b[1],tempResult1[10]);
_2_1_mux_v2 mux_layer1_12(tempResult0[11],tempResult0[13],b[1],tempResult1[11]);
_2_1_mux_v2 mux_layer1_13(tempResult0[12],tempResult0[14],b[1],tempResult1[12]);
_2_1_mux_v2 mux_layer1_14(tempResult0[13],tempResult0[15],b[1],tempResult1[13]);
_2_1_mux_v2 mux_layer1_15(tempResult0[14],tempResult0[16],b[1],tempResult1[14]);
_2_1_mux_v2 mux_layer1_16(tempResult0[15],tempResult0[17],b[1],tempResult1[15]);
_2_1_mux_v2 mux_layer1_17(tempResult0[16],tempResult0[18],b[1],tempResult1[16]);
_2_1_mux_v2 mux_layer1_18(tempResult0[17],tempResult0[19],b[1],tempResult1[17]);
_2_1_mux_v2 mux_layer1_19(tempResult0[18],tempResult0[20],b[1],tempResult1[18]);
_2_1_mux_v2 mux_layer1_20(tempResult0[19],tempResult0[21],b[1],tempResult1[19]);
_2_1_mux_v2 mux_layer1_21(tempResult0[20],tempResult0[22],b[1],tempResult1[20]);
_2_1_mux_v2 mux_layer1_22(tempResult0[21],tempResult0[23],b[1],tempResult1[21]);
_2_1_mux_v2 mux_layer1_23(tempResult0[22],tempResult0[24],b[1],tempResult1[22]);
_2_1_mux_v2 mux_layer1_24(tempResult0[23],tempResult0[25],b[1],tempResult1[23]);
_2_1_mux_v2 mux_layer1_25(tempResult0[24],tempResult0[26],b[1],tempResult1[24]);
_2_1_mux_v2 mux_layer1_26(tempResult0[25],tempResult0[27],b[1],tempResult1[25]);
_2_1_mux_v2 mux_layer1_27(tempResult0[26],tempResult0[28],b[1],tempResult1[26]);
_2_1_mux_v2 mux_layer1_28(tempResult0[27],tempResult0[29],b[1],tempResult1[27]);
_2_1_mux_v2 mux_layer1_29(tempResult0[28],tempResult0[30],b[1],tempResult1[28]);
_2_1_mux_v2 mux_layer1_30(tempResult0[29],tempResult0[31],b[1],tempResult1[29]);
_2_1_mux_v2 mux_layer1_31(tempResult0[30],1'b0,b[1],tempResult1[30]);
_2_1_mux_v2 mux_layer1_32(tempResult0[31],1'b0,b[1],tempResult1[31]);

_2_1_mux_v2 mux_layer2_1(tempResult1[0],tempResult1[4],b[2],tempResult2[0]);
_2_1_mux_v2 mux_layer2_2(tempResult1[1],tempResult1[5],b[2],tempResult2[1]);
_2_1_mux_v2 mux_layer2_3(tempResult1[2],tempResult1[6],b[2],tempResult2[2]);
_2_1_mux_v2 mux_layer2_4(tempResult1[3],tempResult1[7],b[2],tempResult2[3]);
_2_1_mux_v2 mux_layer2_5(tempResult1[4],tempResult1[8],b[2],tempResult2[4]);
_2_1_mux_v2 mux_layer2_6(tempResult1[5],tempResult1[9],b[2],tempResult2[5]);
_2_1_mux_v2 mux_layer2_7(tempResult1[6],tempResult1[10],b[2],tempResult2[6]);
_2_1_mux_v2 mux_layer2_8(tempResult1[7],tempResult1[11],b[2],tempResult2[7]);
_2_1_mux_v2 mux_layer2_9(tempResult1[8],tempResult1[12],b[2],tempResult2[8]);
_2_1_mux_v2 mux_layer2_10(tempResult1[9],tempResult1[13],b[2],tempResult2[9]);
_2_1_mux_v2 mux_layer2_11(tempResult1[10],tempResult1[14],b[2],tempResult2[10]);
_2_1_mux_v2 mux_layer2_12(tempResult1[11],tempResult1[15],b[2],tempResult2[11]);
_2_1_mux_v2 mux_layer2_13(tempResult1[12],tempResult1[16],b[2],tempResult2[12]);
_2_1_mux_v2 mux_layer2_14(tempResult1[13],tempResult1[17],b[2],tempResult2[13]);
_2_1_mux_v2 mux_layer2_15(tempResult1[14],tempResult1[18],b[2],tempResult2[14]);
_2_1_mux_v2 mux_layer2_16(tempResult1[15],tempResult1[19],b[2],tempResult2[15]);
_2_1_mux_v2 mux_layer2_17(tempResult1[16],tempResult1[20],b[2],tempResult2[16]);
_2_1_mux_v2 mux_layer2_18(tempResult1[17],tempResult1[21],b[2],tempResult2[17]);
_2_1_mux_v2 mux_layer2_19(tempResult1[18],tempResult1[22],b[2],tempResult2[18]);
_2_1_mux_v2 mux_layer2_20(tempResult1[19],tempResult1[23],b[2],tempResult2[19]);
_2_1_mux_v2 mux_layer2_21(tempResult1[20],tempResult1[24],b[2],tempResult2[20]);
_2_1_mux_v2 mux_layer2_22(tempResult1[21],tempResult1[25],b[2],tempResult2[21]);
_2_1_mux_v2 mux_layer2_23(tempResult1[22],tempResult1[26],b[2],tempResult2[22]);
_2_1_mux_v2 mux_layer2_24(tempResult1[23],tempResult1[27],b[2],tempResult2[23]);
_2_1_mux_v2 mux_layer2_25(tempResult1[24],tempResult1[28],b[2],tempResult2[24]);
_2_1_mux_v2 mux_layer2_26(tempResult1[25],tempResult1[29],b[2],tempResult2[25]);
_2_1_mux_v2 mux_layer2_27(tempResult1[26],tempResult1[30],b[2],tempResult2[26]);
_2_1_mux_v2 mux_layer2_28(tempResult1[27],tempResult1[31],b[2],tempResult2[27]);
_2_1_mux_v2 mux_layer2_29(tempResult1[28],1'b0,b[2],tempResult2[28]);
_2_1_mux_v2 mux_layer2_30(tempResult1[29],1'b0,b[2],tempResult2[29]);
_2_1_mux_v2 mux_layer2_31(tempResult1[30],1'b0,b[2],tempResult2[30]);
_2_1_mux_v2 mux_layer2_32(tempResult1[31],1'b0,b[2],tempResult2[31]);


_2_1_mux_v2 mux_layer_3_1(tempResult2[0],tempResult2[8],b[3],tempResult3[0]);
_2_1_mux_v2 mux_layer_3_2(tempResult2[1],tempResult2[9],b[3],tempResult3[1]);
_2_1_mux_v2 mux_layer_3_3(tempResult2[2],tempResult2[10],b[3],tempResult3[2]);
_2_1_mux_v2 mux_layer_3_4(tempResult2[3],tempResult2[11],b[3],tempResult3[3]);
_2_1_mux_v2 mux_layer_3_5(tempResult2[4],tempResult2[12],b[3],tempResult3[4]);
_2_1_mux_v2 mux_layer_3_6(tempResult2[5],tempResult2[13],b[3],tempResult3[5]);
_2_1_mux_v2 mux_layer_3_7(tempResult2[6],tempResult2[14],b[3],tempResult3[6]);
_2_1_mux_v2 mux_layer_3_8(tempResult2[7],tempResult2[15],b[3],tempResult3[7]);
_2_1_mux_v2 mux_layer_3_9(tempResult2[8],tempResult2[16],b[3],tempResult3[8]);
_2_1_mux_v2 mux_layer_3_10(tempResult2[9],tempResult2[17],b[3],tempResult3[9]);
_2_1_mux_v2 mux_layer_3_11(tempResult2[10],tempResult2[18],b[3],tempResult3[10]);
_2_1_mux_v2 mux_layer_3_12(tempResult2[11],tempResult2[19],b[3],tempResult3[11]);
_2_1_mux_v2 mux_layer_3_13(tempResult2[12],tempResult2[20],b[3],tempResult3[12]);
_2_1_mux_v2 mux_layer_3_14(tempResult2[13],tempResult2[21],b[3],tempResult3[13]);
_2_1_mux_v2 mux_layer_3_15(tempResult2[14],tempResult2[22],b[3],tempResult3[14]);
_2_1_mux_v2 mux_layer_3_16(tempResult2[15],tempResult2[23],b[3],tempResult3[15]);
_2_1_mux_v2 mux_layer_3_17(tempResult2[16],tempResult2[24],b[3],tempResult3[16]);
_2_1_mux_v2 mux_layer_3_18(tempResult2[17],tempResult2[25],b[3],tempResult3[17]);
_2_1_mux_v2 mux_layer_3_19(tempResult2[18],tempResult2[26],b[3],tempResult3[18]);
_2_1_mux_v2 mux_layer_3_20(tempResult2[19],tempResult2[27],b[3],tempResult3[19]);
_2_1_mux_v2 mux_layer_3_21(tempResult2[20],tempResult2[28],b[3],tempResult3[20]);
_2_1_mux_v2 mux_layer_3_22(tempResult2[21],tempResult2[29],b[3],tempResult3[21]);
_2_1_mux_v2 mux_layer_3_23(tempResult2[22],tempResult2[30],b[3],tempResult3[22]);
_2_1_mux_v2 mux_layer_3_24(tempResult2[23],tempResult2[31],b[3],tempResult3[23]);
_2_1_mux_v2 mux_layer_3_25(tempResult2[24],1'b0,b[3],tempResult3[24]);
_2_1_mux_v2 mux_layer_3_26(tempResult2[25],1'b0,b[3],tempResult3[25]);
_2_1_mux_v2 mux_layer_3_27(tempResult2[26],1'b0,b[3],tempResult3[26]);
_2_1_mux_v2 mux_layer_3_28(tempResult2[27],1'b0,b[3],tempResult3[27]);
_2_1_mux_v2 mux_layer_3_29(tempResult2[28],1'b0,b[3],tempResult3[28]);
_2_1_mux_v2 mux_layer_3_30(tempResult2[29],1'b0,b[3],tempResult3[29]);
_2_1_mux_v2 mux_layer_3_31(tempResult2[30],1'b0,b[3],tempResult3[30]);
_2_1_mux_v2 mux_layer_3_32(tempResult2[31],1'b0,b[3],tempResult3[31]);


_2_1_mux_v2 mux_layer4_1(tempResult3[0],tempResult3[16],b[4],temp_out[0]);
_2_1_mux_v2 mux_layer4_2(tempResult3[1],tempResult3[17],b[4],temp_out[1]);
_2_1_mux_v2 mux_layer4_3(tempResult3[2],tempResult3[18],b[4],temp_out[2]);
_2_1_mux_v2 mux_layer4_4(tempResult3[3],tempResult3[19],b[4],temp_out[3]);
_2_1_mux_v2 mux_layer4_5(tempResult3[4],tempResult3[20],b[4],temp_out[4]);
_2_1_mux_v2 mux_layer4_6(tempResult3[5],tempResult3[21],b[4],temp_out[5]);
_2_1_mux_v2 mux_layer4_7(tempResult3[6],tempResult3[22],b[4],temp_out[6]);
_2_1_mux_v2 mux_layer4_8(tempResult3[7],tempResult3[23],b[4],temp_out[7]);
_2_1_mux_v2 mux_layer4_9(tempResult3[8],tempResult3[24],b[4],temp_out[8]);
_2_1_mux_v2 mux_layer4_10(tempResult3[9],tempResult3[25],b[4],temp_out[9]);
_2_1_mux_v2 mux_layer4_11(tempResult3[10],tempResult3[26],b[4],temp_out[10]);
_2_1_mux_v2 mux_layer4_12(tempResult3[11],tempResult3[27],b[4],temp_out[11]);
_2_1_mux_v2 mux_layer4_13(tempResult3[12],tempResult3[28],b[4],temp_out[12]);
_2_1_mux_v2 mux_layer4_14(tempResult3[13],tempResult3[29],b[4],temp_out[13]);
_2_1_mux_v2 mux_layer4_15(tempResult3[14],tempResult3[30],b[4],temp_out[14]);
_2_1_mux_v2 mux_layer4_16(tempResult3[15],tempResult3[31],b[4],temp_out[15]);
_2_1_mux_v2 mux_layer4_17(tempResult3[16],1'b0,b[4],temp_out[16]);
_2_1_mux_v2 mux_layer4_18(tempResult3[17],1'b0,b[4],temp_out[17]);
_2_1_mux_v2 mux_layer4_19(tempResult3[18],1'b0,b[4],temp_out[18]);
_2_1_mux_v2 mux_layer4_20(tempResult3[19],1'b0,b[4],temp_out[19]);
_2_1_mux_v2 mux_layer4_21(tempResult3[20],1'b0,b[4],temp_out[20]);
_2_1_mux_v2 mux_layer4_22(tempResult3[21],1'b0,b[4],temp_out[21]);
_2_1_mux_v2 mux_layer4_23(tempResult3[22],1'b0,b[4],temp_out[22]);
_2_1_mux_v2 mux_layer4_24(tempResult3[23],1'b0,b[4],temp_out[23]);
_2_1_mux_v2 mux_layer4_25(tempResult3[24],1'b0,b[4],temp_out[24]);
_2_1_mux_v2 mux_layer4_26(tempResult3[25],1'b0,b[4],temp_out[25]);
_2_1_mux_v2 mux_layer4_27(tempResult3[26],1'b0,b[4],temp_out[26]);
_2_1_mux_v2 mux_layer4_28(tempResult3[27],1'b0,b[4],temp_out[27]);
_2_1_mux_v2 mux_layer4_29(tempResult3[28],1'b0,b[4],temp_out[28]);
_2_1_mux_v2 mux_layer4_30(tempResult3[29],1'b0,b[4],temp_out[29]);
_2_1_mux_v2 mux_layer4_31(tempResult3[30],1'b0,b[4],temp_out[30]);
_2_1_mux_v2 mux_layer4_32(tempResult3[31],1'b0,b[4],temp_out[31]);

or or1(overflow,b[5],b[6],b[7],b[8],b[9],b[10],b[11],b[12],b[13],b[14],b[15],b[16],b[17],b[18],b[19],b[20],b[21],b[22],b[23],b[24],b[25],b[26],b[27],b[28],b[29],b[30],b[31]);

not not1(not_overflow,overflow);

and aand0 (out[0],temp_out[0],not_overflow);
and aand1 (out[1],temp_out[1],not_overflow);
and aand2 (out[2],temp_out[2],not_overflow);
and aand3 (out[3],temp_out[3],not_overflow);
and aand4 (out[4],temp_out[4],not_overflow);
and aand5 (out[5],temp_out[5],not_overflow);
and aand6 (out[6],temp_out[6],not_overflow);
and aand7 (out[7],temp_out[7],not_overflow);
and aand8 (out[8],temp_out[8],not_overflow);
and aand9 (out[9],temp_out[9],not_overflow);
and aand10 (out[10],temp_out[10],not_overflow);
and aand11 (out[11],temp_out[11],not_overflow);
and aand12 (out[12],temp_out[12],not_overflow);
and aand13 (out[13],temp_out[13],not_overflow);
and aand14 (out[14],temp_out[14],not_overflow);
and aand15 (out[15],temp_out[15],not_overflow);
and aand16 (out[16],temp_out[16],not_overflow);
and aand17 (out[17],temp_out[17],not_overflow);
and aand18 (out[18],temp_out[18],not_overflow);
and aand19 (out[19],temp_out[19],not_overflow);
and aand20 (out[20],temp_out[20],not_overflow);
and aand21 (out[21],temp_out[21],not_overflow);
and aand22 (out[22],temp_out[22],not_overflow);
and aand23 (out[23],temp_out[23],not_overflow);
and aand24 (out[24],temp_out[24],not_overflow);
and aand25 (out[25],temp_out[25],not_overflow);
and aand26 (out[26],temp_out[26],not_overflow);
and aand27 (out[27],temp_out[27],not_overflow);
and aand28 (out[28],temp_out[28],not_overflow);
and aand29 (out[29],temp_out[29],not_overflow);
and aand30 (out[30],temp_out[30],not_overflow);
and aand31 (out[31],temp_out[31],not_overflow);

endmodule
